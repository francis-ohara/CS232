-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- PROGRAM		"Quartus II 32-bit"
-- VERSION		"Version 13.1.0 Build 162 10/23/2013 SJ Web Edition"
-- CREATED		"Wed Feb 26 20:29:57 2025"

LIBRARY ieee;
USE ieee.std_logic_1164.all; 

LIBRARY work;

ENTITY prime_extension IS 
	PORT
	(
		A :  IN  STD_LOGIC;
		B :  IN  STD_LOGIC;
		C :  IN  STD_LOGIC;
		D :  IN  STD_LOGIC;
		E :  IN  STD_LOGIC;
		O :  OUT  STD_LOGIC
	);
END prime_extension;

ARCHITECTURE bdf_type OF prime_extension IS 

SIGNAL	SYNTHESIZED_WIRE_37 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_38 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_39 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_40 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_41 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_11 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_12 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_13 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_14 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_15 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_16 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_17 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_18 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_19 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_20 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_21 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_22 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_23 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_42 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_43 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_44 :  STD_LOGIC;


BEGIN 



SYNTHESIZED_WIRE_21 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND D AND SYNTHESIZED_WIRE_40 AND SYNTHESIZED_WIRE_40;


SYNTHESIZED_WIRE_19 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND D AND E AND E;


SYNTHESIZED_WIRE_18 <= C AND A AND B AND D AND E AND E;


SYNTHESIZED_WIRE_38 <= NOT(A);



SYNTHESIZED_WIRE_39 <= NOT(B);



SYNTHESIZED_WIRE_37 <= NOT(C);



SYNTHESIZED_WIRE_41 <= NOT(D);



SYNTHESIZED_WIRE_40 <= NOT(E);



SYNTHESIZED_WIRE_43 <= NOT(B);



SYNTHESIZED_WIRE_42 <= NOT(C);



SYNTHESIZED_WIRE_44 <= NOT(D);



SYNTHESIZED_WIRE_20 <= C AND SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND SYNTHESIZED_WIRE_41 AND E AND E;


SYNTHESIZED_WIRE_22 <= SYNTHESIZED_WIRE_11 OR SYNTHESIZED_WIRE_12 OR SYNTHESIZED_WIRE_13 OR SYNTHESIZED_WIRE_14 OR SYNTHESIZED_WIRE_15 OR SYNTHESIZED_WIRE_16 OR SYNTHESIZED_WIRE_17 OR SYNTHESIZED_WIRE_18;


SYNTHESIZED_WIRE_23 <= SYNTHESIZED_WIRE_19 OR SYNTHESIZED_WIRE_20 OR SYNTHESIZED_WIRE_21;


O <= SYNTHESIZED_WIRE_22 OR SYNTHESIZED_WIRE_23;


SYNTHESIZED_WIRE_11 <= C AND SYNTHESIZED_WIRE_38 AND SYNTHESIZED_WIRE_39 AND D AND E AND E;


SYNTHESIZED_WIRE_13 <= SYNTHESIZED_WIRE_37 AND SYNTHESIZED_WIRE_38 AND B AND D AND E AND E;


SYNTHESIZED_WIRE_12 <= C AND SYNTHESIZED_WIRE_38 AND B AND SYNTHESIZED_WIRE_41 AND E AND E;


SYNTHESIZED_WIRE_14 <= SYNTHESIZED_WIRE_42 AND A AND SYNTHESIZED_WIRE_43 AND SYNTHESIZED_WIRE_44 AND E AND E;


SYNTHESIZED_WIRE_16 <= SYNTHESIZED_WIRE_42 AND A AND SYNTHESIZED_WIRE_43 AND D AND E AND E;


SYNTHESIZED_WIRE_15 <= C AND A AND SYNTHESIZED_WIRE_43 AND D AND E AND E;


SYNTHESIZED_WIRE_17 <= C AND A AND B AND SYNTHESIZED_WIRE_44 AND E AND E;


END bdf_type;